// Eric Yeats / Brady Taylor
// ECE 552 Advanced Computer Architecture I
// Final Project
// Fire Fifo


// This module will store the tags of neurons
// that fire in a given time step. The tags are
// stored for processing by the synaptic update proc.

module fire_fifo(
    input clk, 
);
